module();

//this is an empty module
wire a;
wire b = a*2;


endmodule