module();

//this is an empty module

endmodule